module reliability_LUT(
    input   [1:0]   N_channel,
    input   [8:0]   channel_index,
    output  [8:0]   reliability_index
);

    // N = 128 --> 00 10000000
    // N = 256 --> 01 00000000
    // N = 512 --> 10 00000000

    wire [6:0] rindex_128 [0:127];
    wire [7:0] rindex_256 [0:255];
    wire [8:0] rindex_512 [0:511];

    assign reliability_index = (N_channel == 2'b00) ? rindex_128[channel_index] :
                               (N_channel == 2'b01) ? rindex_256[channel_index] :
                                                      rindex_512[channel_index];

    // ===========================================
    //                  N = 128
    // ===========================================

    assign  rindex_128[0] = 0;
    assign  rindex_128[1] = 1;
    assign  rindex_128[2] = 2;
    assign  rindex_128[3] = 4;
    assign  rindex_128[4] = 8;
    assign  rindex_128[5] = 16;
    assign  rindex_128[6] = 32;
    assign  rindex_128[7] = 3;
    assign  rindex_128[8] = 5;
    assign  rindex_128[9] = 64;
    assign  rindex_128[10] = 9;
    assign  rindex_128[11] = 6;
    assign  rindex_128[12] = 17;
    assign  rindex_128[13] = 10;
    assign  rindex_128[14] = 18;
    assign  rindex_128[15] = 12;
    assign  rindex_128[16] = 33;
    assign  rindex_128[17] = 65;
    assign  rindex_128[18] = 20;
    assign  rindex_128[19] = 34;
    assign  rindex_128[20] = 24;
    assign  rindex_128[21] = 36;
    assign  rindex_128[22] = 7;
    assign  rindex_128[23] = 66;
    assign  rindex_128[24] = 11;
    assign  rindex_128[25] = 40;
    assign  rindex_128[26] = 68;
    assign  rindex_128[27] = 19;
    assign  rindex_128[28] = 13;
    assign  rindex_128[29] = 48;
    assign  rindex_128[30] = 14;
    assign  rindex_128[31] = 72;
    assign  rindex_128[32] = 21;
    assign  rindex_128[33] = 35;
    assign  rindex_128[34] = 26;
    assign  rindex_128[35] = 80;
    assign  rindex_128[36] = 37;
    assign  rindex_128[37] = 25;
    assign  rindex_128[38] = 22;
    assign  rindex_128[39] = 38;
    assign  rindex_128[40] = 96;
    assign  rindex_128[41] = 67;
    assign  rindex_128[42] = 41;
    assign  rindex_128[43] = 28;
    assign  rindex_128[44] = 69;
    assign  rindex_128[45] = 42;
    assign  rindex_128[46] = 49;
    assign  rindex_128[47] = 74;
    assign  rindex_128[48] = 70;
    assign  rindex_128[49] = 44;
    assign  rindex_128[50] = 81;
    assign  rindex_128[51] = 50;
    assign  rindex_128[52] = 73;
    assign  rindex_128[53] = 15;
    assign  rindex_128[54] = 52;
    assign  rindex_128[55] = 23;
    assign  rindex_128[56] = 76;
    assign  rindex_128[57] = 82;
    assign  rindex_128[58] = 56;
    assign  rindex_128[59] = 27;
    assign  rindex_128[60] = 97;
    assign  rindex_128[61] = 39;
    assign  rindex_128[62] = 84;
    assign  rindex_128[63] = 29;
    assign  rindex_128[64] = 43;
    assign  rindex_128[65] = 98;
    assign  rindex_128[66] = 88;
    assign  rindex_128[67] = 30;
    assign  rindex_128[68] = 71;
    assign  rindex_128[69] = 45;
    assign  rindex_128[70] = 100;
    assign  rindex_128[71] = 51;
    assign  rindex_128[72] = 46;
    assign  rindex_128[73] = 75;
    assign  rindex_128[74] = 104;
    assign  rindex_128[75] = 53;
    assign  rindex_128[76] = 77;
    assign  rindex_128[77] = 54;
    assign  rindex_128[78] = 83;
    assign  rindex_128[79] = 57;
    assign  rindex_128[80] = 112;
    assign  rindex_128[81] = 78;
    assign  rindex_128[82] = 85;
    assign  rindex_128[83] = 58;
    assign  rindex_128[84] = 99;
    assign  rindex_128[85] = 86;
    assign  rindex_128[86] = 60;
    assign  rindex_128[87] = 89;
    assign  rindex_128[88] = 101;
    assign  rindex_128[89] = 31;
    assign  rindex_128[90] = 90;
    assign  rindex_128[91] = 102;
    assign  rindex_128[92] = 105;
    assign  rindex_128[93] = 92;
    assign  rindex_128[94] = 47;
    assign  rindex_128[95] = 106;
    assign  rindex_128[96] = 55;
    assign  rindex_128[97] = 113;
    assign  rindex_128[98] = 79;
    assign  rindex_128[99] = 108;
    assign  rindex_128[100] = 59;
    assign  rindex_128[101] = 114;
    assign  rindex_128[102] = 87;
    assign  rindex_128[103] = 116;
    assign  rindex_128[104] = 61;
    assign  rindex_128[105] = 91;
    assign  rindex_128[106] = 120;
    assign  rindex_128[107] = 62;
    assign  rindex_128[108] = 103;
    assign  rindex_128[109] = 93;
    assign  rindex_128[110] = 107;
    assign  rindex_128[111] = 94;
    assign  rindex_128[112] = 109;
    assign  rindex_128[113] = 115;
    assign  rindex_128[114] = 110;
    assign  rindex_128[115] = 117;
    assign  rindex_128[116] = 118;
    assign  rindex_128[117] = 121;
    assign  rindex_128[118] = 122;
    assign  rindex_128[119] = 63;
    assign  rindex_128[120] = 124;
    assign  rindex_128[121] = 95;
    assign  rindex_128[122] = 111;
    assign  rindex_128[123] = 119;
    assign  rindex_128[124] = 123;
    assign  rindex_128[125] = 125;
    assign  rindex_128[126] = 126;
    assign  rindex_128[127] = 127;
    
    // ===========================================
    //                  N = 256
    // ===========================================

    assign  rindex_256[0] = 0;
    assign  rindex_256[1] = 1;
    assign  rindex_256[2] = 2;
    assign  rindex_256[3] = 4;
    assign  rindex_256[4] = 8;
    assign  rindex_256[5] = 16;
    assign  rindex_256[6] = 32;
    assign  rindex_256[7] = 3;
    assign  rindex_256[8] = 5;
    assign  rindex_256[9] = 64;
    assign  rindex_256[10] = 9;
    assign  rindex_256[11] = 6;
    assign  rindex_256[12] = 17;
    assign  rindex_256[13] = 10;
    assign  rindex_256[14] = 18;
    assign  rindex_256[15] = 128;
    assign  rindex_256[16] = 12;
    assign  rindex_256[17] = 33;
    assign  rindex_256[18] = 65;
    assign  rindex_256[19] = 20;
    assign  rindex_256[20] = 34;
    assign  rindex_256[21] = 24;
    assign  rindex_256[22] = 36;
    assign  rindex_256[23] = 7;
    assign  rindex_256[24] = 129;
    assign  rindex_256[25] = 66;
    assign  rindex_256[26] = 11;
    assign  rindex_256[27] = 40;
    assign  rindex_256[28] = 68;
    assign  rindex_256[29] = 130;
    assign  rindex_256[30] = 19;
    assign  rindex_256[31] = 13;
    assign  rindex_256[32] = 48;
    assign  rindex_256[33] = 14;
    assign  rindex_256[34] = 72;
    assign  rindex_256[35] = 21;
    assign  rindex_256[36] = 132;
    assign  rindex_256[37] = 35;
    assign  rindex_256[38] = 26;
    assign  rindex_256[39] = 80;
    assign  rindex_256[40] = 37;
    assign  rindex_256[41] = 25;
    assign  rindex_256[42] = 22;
    assign  rindex_256[43] = 136;
    assign  rindex_256[44] = 38;
    assign  rindex_256[45] = 96;
    assign  rindex_256[46] = 67;
    assign  rindex_256[47] = 41;
    assign  rindex_256[48] = 144;
    assign  rindex_256[49] = 28;
    assign  rindex_256[50] = 69;
    assign  rindex_256[51] = 42;
    assign  rindex_256[52] = 49;
    assign  rindex_256[53] = 74;
    assign  rindex_256[54] = 160;
    assign  rindex_256[55] = 192;
    assign  rindex_256[56] = 70;
    assign  rindex_256[57] = 44;
    assign  rindex_256[58] = 131;
    assign  rindex_256[59] = 81;
    assign  rindex_256[60] = 50;
    assign  rindex_256[61] = 73;
    assign  rindex_256[62] = 15;
    assign  rindex_256[63] = 133;
    assign  rindex_256[64] = 52;
    assign  rindex_256[65] = 23;
    assign  rindex_256[66] = 134;
    assign  rindex_256[67] = 76;
    assign  rindex_256[68] = 137;
    assign  rindex_256[69] = 82;
    assign  rindex_256[70] = 56;
    assign  rindex_256[71] = 27;
    assign  rindex_256[72] = 97;
    assign  rindex_256[73] = 39;
    assign  rindex_256[74] = 84;
    assign  rindex_256[75] = 138;
    assign  rindex_256[76] = 145;
    assign  rindex_256[77] = 29;
    assign  rindex_256[78] = 43;
    assign  rindex_256[79] = 98;
    assign  rindex_256[80] = 88;
    assign  rindex_256[81] = 140;
    assign  rindex_256[82] = 30;
    assign  rindex_256[83] = 146;
    assign  rindex_256[84] = 71;
    assign  rindex_256[85] = 161;
    assign  rindex_256[86] = 45;
    assign  rindex_256[87] = 100;
    assign  rindex_256[88] = 51;
    assign  rindex_256[89] = 148;
    assign  rindex_256[90] = 46;
    assign  rindex_256[91] = 75;
    assign  rindex_256[92] = 104;
    assign  rindex_256[93] = 162;
    assign  rindex_256[94] = 53;
    assign  rindex_256[95] = 193;
    assign  rindex_256[96] = 152;
    assign  rindex_256[97] = 77;
    assign  rindex_256[98] = 164;
    assign  rindex_256[99] = 54;
    assign  rindex_256[100] = 83;
    assign  rindex_256[101] = 57;
    assign  rindex_256[102] = 112;
    assign  rindex_256[103] = 135;
    assign  rindex_256[104] = 78;
    assign  rindex_256[105] = 194;
    assign  rindex_256[106] = 85;
    assign  rindex_256[107] = 58;
    assign  rindex_256[108] = 168;
    assign  rindex_256[109] = 139;
    assign  rindex_256[110] = 99;
    assign  rindex_256[111] = 86;
    assign  rindex_256[112] = 60;
    assign  rindex_256[113] = 89;
    assign  rindex_256[114] = 196;
    assign  rindex_256[115] = 141;
    assign  rindex_256[116] = 101;
    assign  rindex_256[117] = 147;
    assign  rindex_256[118] = 176;
    assign  rindex_256[119] = 142;
    assign  rindex_256[120] = 31;
    assign  rindex_256[121] = 200;
    assign  rindex_256[122] = 90;
    assign  rindex_256[123] = 149;
    assign  rindex_256[124] = 102;
    assign  rindex_256[125] = 105;
    assign  rindex_256[126] = 163;
    assign  rindex_256[127] = 92;
    assign  rindex_256[128] = 47;
    assign  rindex_256[129] = 208;
    assign  rindex_256[130] = 150;
    assign  rindex_256[131] = 153;
    assign  rindex_256[132] = 165;
    assign  rindex_256[133] = 106;
    assign  rindex_256[134] = 55;
    assign  rindex_256[135] = 113;
    assign  rindex_256[136] = 154;
    assign  rindex_256[137] = 79;
    assign  rindex_256[138] = 108;
    assign  rindex_256[139] = 224;
    assign  rindex_256[140] = 166;
    assign  rindex_256[141] = 195;
    assign  rindex_256[142] = 59;
    assign  rindex_256[143] = 169;
    assign  rindex_256[144] = 114;
    assign  rindex_256[145] = 156;
    assign  rindex_256[146] = 87;
    assign  rindex_256[147] = 197;
    assign  rindex_256[148] = 116;
    assign  rindex_256[149] = 170;
    assign  rindex_256[150] = 61;
    assign  rindex_256[151] = 177;
    assign  rindex_256[152] = 91;
    assign  rindex_256[153] = 198;
    assign  rindex_256[154] = 172;
    assign  rindex_256[155] = 120;
    assign  rindex_256[156] = 201;
    assign  rindex_256[157] = 62;
    assign  rindex_256[158] = 143;
    assign  rindex_256[159] = 103;
    assign  rindex_256[160] = 178;
    assign  rindex_256[161] = 93;
    assign  rindex_256[162] = 202;
    assign  rindex_256[163] = 107;
    assign  rindex_256[164] = 180;
    assign  rindex_256[165] = 151;
    assign  rindex_256[166] = 209;
    assign  rindex_256[167] = 94;
    assign  rindex_256[168] = 204;
    assign  rindex_256[169] = 155;
    assign  rindex_256[170] = 210;
    assign  rindex_256[171] = 109;
    assign  rindex_256[172] = 184;
    assign  rindex_256[173] = 115;
    assign  rindex_256[174] = 167;
    assign  rindex_256[175] = 225;
    assign  rindex_256[176] = 157;
    assign  rindex_256[177] = 110;
    assign  rindex_256[178] = 117;
    assign  rindex_256[179] = 212;
    assign  rindex_256[180] = 171;
    assign  rindex_256[181] = 226;
    assign  rindex_256[182] = 216;
    assign  rindex_256[183] = 158;
    assign  rindex_256[184] = 118;
    assign  rindex_256[185] = 173;
    assign  rindex_256[186] = 121;
    assign  rindex_256[187] = 199;
    assign  rindex_256[188] = 179;
    assign  rindex_256[189] = 228;
    assign  rindex_256[190] = 174;
    assign  rindex_256[191] = 122;
    assign  rindex_256[192] = 203;
    assign  rindex_256[193] = 63;
    assign  rindex_256[194] = 181;
    assign  rindex_256[195] = 232;
    assign  rindex_256[196] = 124;
    assign  rindex_256[197] = 205;
    assign  rindex_256[198] = 182;
    assign  rindex_256[199] = 211;
    assign  rindex_256[200] = 185;
    assign  rindex_256[201] = 240;
    assign  rindex_256[202] = 206;
    assign  rindex_256[203] = 95;
    assign  rindex_256[204] = 213;
    assign  rindex_256[205] = 186;
    assign  rindex_256[206] = 227;
    assign  rindex_256[207] = 111;
    assign  rindex_256[208] = 214;
    assign  rindex_256[209] = 188;
    assign  rindex_256[210] = 217;
    assign  rindex_256[211] = 229;
    assign  rindex_256[212] = 159;
    assign  rindex_256[213] = 119;
    assign  rindex_256[214] = 218;
    assign  rindex_256[215] = 230;
    assign  rindex_256[216] = 233;
    assign  rindex_256[217] = 175;
    assign  rindex_256[218] = 123;
    assign  rindex_256[219] = 220;
    assign  rindex_256[220] = 183;
    assign  rindex_256[221] = 234;
    assign  rindex_256[222] = 125;
    assign  rindex_256[223] = 241;
    assign  rindex_256[224] = 207;
    assign  rindex_256[225] = 187;
    assign  rindex_256[226] = 236;
    assign  rindex_256[227] = 126;
    assign  rindex_256[228] = 242;
    assign  rindex_256[229] = 244;
    assign  rindex_256[230] = 189;
    assign  rindex_256[231] = 215;
    assign  rindex_256[232] = 219;
    assign  rindex_256[233] = 231;
    assign  rindex_256[234] = 248;
    assign  rindex_256[235] = 190;
    assign  rindex_256[236] = 221;
    assign  rindex_256[237] = 235;
    assign  rindex_256[238] = 222;
    assign  rindex_256[239] = 237;
    assign  rindex_256[240] = 243;
    assign  rindex_256[241] = 238;
    assign  rindex_256[242] = 245;
    assign  rindex_256[243] = 127;
    assign  rindex_256[244] = 191;
    assign  rindex_256[245] = 246;
    assign  rindex_256[246] = 249;
    assign  rindex_256[247] = 250;
    assign  rindex_256[248] = 252;
    assign  rindex_256[249] = 223;
    assign  rindex_256[250] = 239;
    assign  rindex_256[251] = 251;
    assign  rindex_256[252] = 247;
    assign  rindex_256[253] = 253;
    assign  rindex_256[254] = 254;
    assign  rindex_256[255] = 255;

    // ===========================================
    //                  N = 512
    // ===========================================

    assign  rindex_512[0] = 0;
    assign  rindex_512[1] = 1;
    assign  rindex_512[2] = 2;
    assign  rindex_512[3] = 4;
    assign  rindex_512[4] = 8;
    assign  rindex_512[5] = 16;
    assign  rindex_512[6] = 32;
    assign  rindex_512[7] = 3;
    assign  rindex_512[8] = 5;
    assign  rindex_512[9] = 64;
    assign  rindex_512[10] = 9;
    assign  rindex_512[11] = 6;
    assign  rindex_512[12] = 17;
    assign  rindex_512[13] = 10;
    assign  rindex_512[14] = 18;
    assign  rindex_512[15] = 128;
    assign  rindex_512[16] = 12;
    assign  rindex_512[17] = 33;
    assign  rindex_512[18] = 65;
    assign  rindex_512[19] = 20;
    assign  rindex_512[20] = 256;
    assign  rindex_512[21] = 34;
    assign  rindex_512[22] = 24;
    assign  rindex_512[23] = 36;
    assign  rindex_512[24] = 7;
    assign  rindex_512[25] = 129;
    assign  rindex_512[26] = 66;
    assign  rindex_512[27] = 11;
    assign  rindex_512[28] = 40;
    assign  rindex_512[29] = 68;
    assign  rindex_512[30] = 130;
    assign  rindex_512[31] = 19;
    assign  rindex_512[32] = 13;
    assign  rindex_512[33] = 48;
    assign  rindex_512[34] = 14;
    assign  rindex_512[35] = 72;
    assign  rindex_512[36] = 257;
    assign  rindex_512[37] = 21;
    assign  rindex_512[38] = 132;
    assign  rindex_512[39] = 35;
    assign  rindex_512[40] = 258;
    assign  rindex_512[41] = 26;
    assign  rindex_512[42] = 80;
    assign  rindex_512[43] = 37;
    assign  rindex_512[44] = 25;
    assign  rindex_512[45] = 22;
    assign  rindex_512[46] = 136;
    assign  rindex_512[47] = 260;
    assign  rindex_512[48] = 264;
    assign  rindex_512[49] = 38;
    assign  rindex_512[50] = 96;
    assign  rindex_512[51] = 67;
    assign  rindex_512[52] = 41;
    assign  rindex_512[53] = 144;
    assign  rindex_512[54] = 28;
    assign  rindex_512[55] = 69;
    assign  rindex_512[56] = 42;
    assign  rindex_512[57] = 49;
    assign  rindex_512[58] = 74;
    assign  rindex_512[59] = 272;
    assign  rindex_512[60] = 160;
    assign  rindex_512[61] = 288;
    assign  rindex_512[62] = 192;
    assign  rindex_512[63] = 70;
    assign  rindex_512[64] = 44;
    assign  rindex_512[65] = 131;
    assign  rindex_512[66] = 81;
    assign  rindex_512[67] = 50;
    assign  rindex_512[68] = 73;
    assign  rindex_512[69] = 15;
    assign  rindex_512[70] = 320;
    assign  rindex_512[71] = 133;
    assign  rindex_512[72] = 52;
    assign  rindex_512[73] = 23;
    assign  rindex_512[74] = 134;
    assign  rindex_512[75] = 384;
    assign  rindex_512[76] = 76;
    assign  rindex_512[77] = 137;
    assign  rindex_512[78] = 82;
    assign  rindex_512[79] = 56;
    assign  rindex_512[80] = 27;
    assign  rindex_512[81] = 97;
    assign  rindex_512[82] = 39;
    assign  rindex_512[83] = 259;
    assign  rindex_512[84] = 84;
    assign  rindex_512[85] = 138;
    assign  rindex_512[86] = 145;
    assign  rindex_512[87] = 261;
    assign  rindex_512[88] = 29;
    assign  rindex_512[89] = 43;
    assign  rindex_512[90] = 98;
    assign  rindex_512[91] = 88;
    assign  rindex_512[92] = 140;
    assign  rindex_512[93] = 30;
    assign  rindex_512[94] = 146;
    assign  rindex_512[95] = 71;
    assign  rindex_512[96] = 262;
    assign  rindex_512[97] = 265;
    assign  rindex_512[98] = 161;
    assign  rindex_512[99] = 45;
    assign  rindex_512[100] = 100;
    assign  rindex_512[101] = 51;
    assign  rindex_512[102] = 148;
    assign  rindex_512[103] = 46;
    assign  rindex_512[104] = 75;
    assign  rindex_512[105] = 266;
    assign  rindex_512[106] = 273;
    assign  rindex_512[107] = 104;
    assign  rindex_512[108] = 162;
    assign  rindex_512[109] = 53;
    assign  rindex_512[110] = 193;
    assign  rindex_512[111] = 152;
    assign  rindex_512[112] = 77;
    assign  rindex_512[113] = 164;
    assign  rindex_512[114] = 268;
    assign  rindex_512[115] = 274;
    assign  rindex_512[116] = 54;
    assign  rindex_512[117] = 83;
    assign  rindex_512[118] = 57;
    assign  rindex_512[119] = 112;
    assign  rindex_512[120] = 135;
    assign  rindex_512[121] = 78;
    assign  rindex_512[122] = 289;
    assign  rindex_512[123] = 194;
    assign  rindex_512[124] = 85;
    assign  rindex_512[125] = 276;
    assign  rindex_512[126] = 58;
    assign  rindex_512[127] = 168;
    assign  rindex_512[128] = 139;
    assign  rindex_512[129] = 99;
    assign  rindex_512[130] = 86;
    assign  rindex_512[131] = 60;
    assign  rindex_512[132] = 280;
    assign  rindex_512[133] = 89;
    assign  rindex_512[134] = 290;
    assign  rindex_512[135] = 196;
    assign  rindex_512[136] = 141;
    assign  rindex_512[137] = 101;
    assign  rindex_512[138] = 147;
    assign  rindex_512[139] = 176;
    assign  rindex_512[140] = 142;
    assign  rindex_512[141] = 321;
    assign  rindex_512[142] = 31;
    assign  rindex_512[143] = 200;
    assign  rindex_512[144] = 90;
    assign  rindex_512[145] = 292;
    assign  rindex_512[146] = 322;
    assign  rindex_512[147] = 263;
    assign  rindex_512[148] = 149;
    assign  rindex_512[149] = 102;
    assign  rindex_512[150] = 105;
    assign  rindex_512[151] = 304;
    assign  rindex_512[152] = 296;
    assign  rindex_512[153] = 163;
    assign  rindex_512[154] = 92;
    assign  rindex_512[155] = 47;
    assign  rindex_512[156] = 267;
    assign  rindex_512[157] = 385;
    assign  rindex_512[158] = 324;
    assign  rindex_512[159] = 208;
    assign  rindex_512[160] = 386;
    assign  rindex_512[161] = 150;
    assign  rindex_512[162] = 153;
    assign  rindex_512[163] = 165;
    assign  rindex_512[164] = 106;
    assign  rindex_512[165] = 55;
    assign  rindex_512[166] = 328;
    assign  rindex_512[167] = 113;
    assign  rindex_512[168] = 154;
    assign  rindex_512[169] = 79;
    assign  rindex_512[170] = 269;
    assign  rindex_512[171] = 108;
    assign  rindex_512[172] = 224;
    assign  rindex_512[173] = 166;
    assign  rindex_512[174] = 195;
    assign  rindex_512[175] = 270;
    assign  rindex_512[176] = 275;
    assign  rindex_512[177] = 291;
    assign  rindex_512[178] = 59;
    assign  rindex_512[179] = 169;
    assign  rindex_512[180] = 114;
    assign  rindex_512[181] = 277;
    assign  rindex_512[182] = 156;
    assign  rindex_512[183] = 87;
    assign  rindex_512[184] = 197;
    assign  rindex_512[185] = 116;
    assign  rindex_512[186] = 170;
    assign  rindex_512[187] = 61;
    assign  rindex_512[188] = 281;
    assign  rindex_512[189] = 278;
    assign  rindex_512[190] = 177;
    assign  rindex_512[191] = 293;
    assign  rindex_512[192] = 388;
    assign  rindex_512[193] = 91;
    assign  rindex_512[194] = 198;
    assign  rindex_512[195] = 172;
    assign  rindex_512[196] = 120;
    assign  rindex_512[197] = 201;
    assign  rindex_512[198] = 336;
    assign  rindex_512[199] = 62;
    assign  rindex_512[200] = 282;
    assign  rindex_512[201] = 143;
    assign  rindex_512[202] = 103;
    assign  rindex_512[203] = 178;
    assign  rindex_512[204] = 294;
    assign  rindex_512[205] = 93;
    assign  rindex_512[206] = 202;
    assign  rindex_512[207] = 323;
    assign  rindex_512[208] = 392;
    assign  rindex_512[209] = 297;
    assign  rindex_512[210] = 107;
    assign  rindex_512[211] = 180;
    assign  rindex_512[212] = 151;
    assign  rindex_512[213] = 209;
    assign  rindex_512[214] = 284;
    assign  rindex_512[215] = 94;
    assign  rindex_512[216] = 204;
    assign  rindex_512[217] = 298;
    assign  rindex_512[218] = 400;
    assign  rindex_512[219] = 352;
    assign  rindex_512[220] = 325;
    assign  rindex_512[221] = 155;
    assign  rindex_512[222] = 210;
    assign  rindex_512[223] = 305;
    assign  rindex_512[224] = 300;
    assign  rindex_512[225] = 109;
    assign  rindex_512[226] = 184;
    assign  rindex_512[227] = 115;
    assign  rindex_512[228] = 167;
    assign  rindex_512[229] = 225;
    assign  rindex_512[230] = 326;
    assign  rindex_512[231] = 306;
    assign  rindex_512[232] = 157;
    assign  rindex_512[233] = 329;
    assign  rindex_512[234] = 110;
    assign  rindex_512[235] = 117;
    assign  rindex_512[236] = 212;
    assign  rindex_512[237] = 171;
    assign  rindex_512[238] = 330;
    assign  rindex_512[239] = 226;
    assign  rindex_512[240] = 387;
    assign  rindex_512[241] = 308;
    assign  rindex_512[242] = 216;
    assign  rindex_512[243] = 416;
    assign  rindex_512[244] = 271;
    assign  rindex_512[245] = 279;
    assign  rindex_512[246] = 158;
    assign  rindex_512[247] = 337;
    assign  rindex_512[248] = 118;
    assign  rindex_512[249] = 332;
    assign  rindex_512[250] = 389;
    assign  rindex_512[251] = 173;
    assign  rindex_512[252] = 121;
    assign  rindex_512[253] = 199;
    assign  rindex_512[254] = 179;
    assign  rindex_512[255] = 228;
    assign  rindex_512[256] = 338;
    assign  rindex_512[257] = 312;
    assign  rindex_512[258] = 390;
    assign  rindex_512[259] = 174;
    assign  rindex_512[260] = 393;
    assign  rindex_512[261] = 283;
    assign  rindex_512[262] = 122;
    assign  rindex_512[263] = 448;
    assign  rindex_512[264] = 353;
    assign  rindex_512[265] = 203;
    assign  rindex_512[266] = 63;
    assign  rindex_512[267] = 340;
    assign  rindex_512[268] = 394;
    assign  rindex_512[269] = 181;
    assign  rindex_512[270] = 295;
    assign  rindex_512[271] = 285;
    assign  rindex_512[272] = 232;
    assign  rindex_512[273] = 124;
    assign  rindex_512[274] = 205;
    assign  rindex_512[275] = 182;
    assign  rindex_512[276] = 286;
    assign  rindex_512[277] = 299;
    assign  rindex_512[278] = 354;
    assign  rindex_512[279] = 211;
    assign  rindex_512[280] = 401;
    assign  rindex_512[281] = 185;
    assign  rindex_512[282] = 396;
    assign  rindex_512[283] = 344;
    assign  rindex_512[284] = 240;
    assign  rindex_512[285] = 206;
    assign  rindex_512[286] = 95;
    assign  rindex_512[287] = 327;
    assign  rindex_512[288] = 402;
    assign  rindex_512[289] = 356;
    assign  rindex_512[290] = 307;
    assign  rindex_512[291] = 301;
    assign  rindex_512[292] = 417;
    assign  rindex_512[293] = 213;
    assign  rindex_512[294] = 186;
    assign  rindex_512[295] = 404;
    assign  rindex_512[296] = 227;
    assign  rindex_512[297] = 418;
    assign  rindex_512[298] = 302;
    assign  rindex_512[299] = 360;
    assign  rindex_512[300] = 111;
    assign  rindex_512[301] = 331;
    assign  rindex_512[302] = 214;
    assign  rindex_512[303] = 309;
    assign  rindex_512[304] = 188;
    assign  rindex_512[305] = 449;
    assign  rindex_512[306] = 217;
    assign  rindex_512[307] = 408;
    assign  rindex_512[308] = 229;
    assign  rindex_512[309] = 159;
    assign  rindex_512[310] = 420;
    assign  rindex_512[311] = 310;
    assign  rindex_512[312] = 333;
    assign  rindex_512[313] = 119;
    assign  rindex_512[314] = 339;
    assign  rindex_512[315] = 218;
    assign  rindex_512[316] = 368;
    assign  rindex_512[317] = 230;
    assign  rindex_512[318] = 391;
    assign  rindex_512[319] = 313;
    assign  rindex_512[320] = 450;
    assign  rindex_512[321] = 334;
    assign  rindex_512[322] = 233;
    assign  rindex_512[323] = 175;
    assign  rindex_512[324] = 123;
    assign  rindex_512[325] = 341;
    assign  rindex_512[326] = 220;
    assign  rindex_512[327] = 314;
    assign  rindex_512[328] = 424;
    assign  rindex_512[329] = 395;
    assign  rindex_512[330] = 355;
    assign  rindex_512[331] = 287;
    assign  rindex_512[332] = 183;
    assign  rindex_512[333] = 234;
    assign  rindex_512[334] = 125;
    assign  rindex_512[335] = 342;
    assign  rindex_512[336] = 316;
    assign  rindex_512[337] = 241;
    assign  rindex_512[338] = 345;
    assign  rindex_512[339] = 452;
    assign  rindex_512[340] = 397;
    assign  rindex_512[341] = 403;
    assign  rindex_512[342] = 207;
    assign  rindex_512[343] = 432;
    assign  rindex_512[344] = 357;
    assign  rindex_512[345] = 187;
    assign  rindex_512[346] = 236;
    assign  rindex_512[347] = 126;
    assign  rindex_512[348] = 242;
    assign  rindex_512[349] = 398;
    assign  rindex_512[350] = 346;
    assign  rindex_512[351] = 456;
    assign  rindex_512[352] = 358;
    assign  rindex_512[353] = 405;
    assign  rindex_512[354] = 303;
    assign  rindex_512[355] = 244;
    assign  rindex_512[356] = 189;
    assign  rindex_512[357] = 361;
    assign  rindex_512[358] = 215;
    assign  rindex_512[359] = 348;
    assign  rindex_512[360] = 419;
    assign  rindex_512[361] = 406;
    assign  rindex_512[362] = 464;
    assign  rindex_512[363] = 362;
    assign  rindex_512[364] = 409;
    assign  rindex_512[365] = 219;
    assign  rindex_512[366] = 311;
    assign  rindex_512[367] = 421;
    assign  rindex_512[368] = 410;
    assign  rindex_512[369] = 231;
    assign  rindex_512[370] = 248;
    assign  rindex_512[371] = 369;
    assign  rindex_512[372] = 190;
    assign  rindex_512[373] = 364;
    assign  rindex_512[374] = 335;
    assign  rindex_512[375] = 480;
    assign  rindex_512[376] = 315;
    assign  rindex_512[377] = 221;
    assign  rindex_512[378] = 370;
    assign  rindex_512[379] = 422;
    assign  rindex_512[380] = 425;
    assign  rindex_512[381] = 451;
    assign  rindex_512[382] = 235;
    assign  rindex_512[383] = 412;
    assign  rindex_512[384] = 343;
    assign  rindex_512[385] = 372;
    assign  rindex_512[386] = 317;
    assign  rindex_512[387] = 222;
    assign  rindex_512[388] = 426;
    assign  rindex_512[389] = 453;
    assign  rindex_512[390] = 237;
    assign  rindex_512[391] = 433;
    assign  rindex_512[392] = 347;
    assign  rindex_512[393] = 243;
    assign  rindex_512[394] = 454;
    assign  rindex_512[395] = 318;
    assign  rindex_512[396] = 376;
    assign  rindex_512[397] = 428;
    assign  rindex_512[398] = 238;
    assign  rindex_512[399] = 359;
    assign  rindex_512[400] = 457;
    assign  rindex_512[401] = 399;
    assign  rindex_512[402] = 434;
    assign  rindex_512[403] = 349;
    assign  rindex_512[404] = 245;
    assign  rindex_512[405] = 458;
    assign  rindex_512[406] = 363;
    assign  rindex_512[407] = 127;
    assign  rindex_512[408] = 191;
    assign  rindex_512[409] = 407;
    assign  rindex_512[410] = 436;
    assign  rindex_512[411] = 465;
    assign  rindex_512[412] = 246;
    assign  rindex_512[413] = 350;
    assign  rindex_512[414] = 460;
    assign  rindex_512[415] = 249;
    assign  rindex_512[416] = 411;
    assign  rindex_512[417] = 365;
    assign  rindex_512[418] = 440;
    assign  rindex_512[419] = 374;
    assign  rindex_512[420] = 423;
    assign  rindex_512[421] = 466;
    assign  rindex_512[422] = 250;
    assign  rindex_512[423] = 371;
    assign  rindex_512[424] = 481;
    assign  rindex_512[425] = 413;
    assign  rindex_512[426] = 366;
    assign  rindex_512[427] = 468;
    assign  rindex_512[428] = 429;
    assign  rindex_512[429] = 252;
    assign  rindex_512[430] = 373;
    assign  rindex_512[431] = 482;
    assign  rindex_512[432] = 427;
    assign  rindex_512[433] = 414;
    assign  rindex_512[434] = 223;
    assign  rindex_512[435] = 472;
    assign  rindex_512[436] = 455;
    assign  rindex_512[437] = 377;
    assign  rindex_512[438] = 435;
    assign  rindex_512[439] = 319;
    assign  rindex_512[440] = 484;
    assign  rindex_512[441] = 430;
    assign  rindex_512[442] = 488;
    assign  rindex_512[443] = 239;
    assign  rindex_512[444] = 378;
    assign  rindex_512[445] = 459;
    assign  rindex_512[446] = 437;
    assign  rindex_512[447] = 380;
    assign  rindex_512[448] = 461;
    assign  rindex_512[449] = 496;
    assign  rindex_512[450] = 351;
    assign  rindex_512[451] = 467;
    assign  rindex_512[452] = 438;
    assign  rindex_512[453] = 251;
    assign  rindex_512[454] = 462;
    assign  rindex_512[455] = 442;
    assign  rindex_512[456] = 441;
    assign  rindex_512[457] = 469;
    assign  rindex_512[458] = 247;
    assign  rindex_512[459] = 367;
    assign  rindex_512[460] = 253;
    assign  rindex_512[461] = 375;
    assign  rindex_512[462] = 444;
    assign  rindex_512[463] = 470;
    assign  rindex_512[464] = 483;
    assign  rindex_512[465] = 415;
    assign  rindex_512[466] = 485;
    assign  rindex_512[467] = 473;
    assign  rindex_512[468] = 474;
    assign  rindex_512[469] = 254;
    assign  rindex_512[470] = 379;
    assign  rindex_512[471] = 431;
    assign  rindex_512[472] = 489;
    assign  rindex_512[473] = 486;
    assign  rindex_512[474] = 476;
    assign  rindex_512[475] = 439;
    assign  rindex_512[476] = 490;
    assign  rindex_512[477] = 463;
    assign  rindex_512[478] = 381;
    assign  rindex_512[479] = 497;
    assign  rindex_512[480] = 492;
    assign  rindex_512[481] = 443;
    assign  rindex_512[482] = 382;
    assign  rindex_512[483] = 498;
    assign  rindex_512[484] = 445;
    assign  rindex_512[485] = 471;
    assign  rindex_512[486] = 500;
    assign  rindex_512[487] = 446;
    assign  rindex_512[488] = 475;
    assign  rindex_512[489] = 487;
    assign  rindex_512[490] = 504;
    assign  rindex_512[491] = 255;
    assign  rindex_512[492] = 477;
    assign  rindex_512[493] = 491;
    assign  rindex_512[494] = 478;
    assign  rindex_512[495] = 383;
    assign  rindex_512[496] = 493;
    assign  rindex_512[497] = 499;
    assign  rindex_512[498] = 502;
    assign  rindex_512[499] = 494;
    assign  rindex_512[500] = 501;
    assign  rindex_512[501] = 447;
    assign  rindex_512[502] = 505;
    assign  rindex_512[503] = 506;
    assign  rindex_512[504] = 479;
    assign  rindex_512[505] = 508;
    assign  rindex_512[506] = 495;
    assign  rindex_512[507] = 503;
    assign  rindex_512[508] = 507;
    assign  rindex_512[509] = 509;
    assign  rindex_512[510] = 510;
    assign  rindex_512[511] = 511;

endmodule
